library verilog;
use verilog.vl_types.all;
entity mem_test_vtf is
end mem_test_vtf;
