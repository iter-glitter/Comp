`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   19:09:37 02/18/2013
// Design Name:   ld_st_shift_nbit
// Module Name:   D:/Users/Hendren/My Documents/School/EE480/DVHW7/ld_st_shift_nbit/ld_st_shift_nbit_vtf.v
// Project Name:  ld_st_shift_nbit
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: ld_st_shift_nbit
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module ld_st_shift_nbit_vtf;

	// Inputs
	reg clk;
	reg clr;
	reg set;
	reg [1:0] ctrl;
	reg ls;
	reg rs;
	reg [3:0] reg_in;
	
	// Outputs
	wire [3:0] reg_out;
	reg [3:0] reg_out_tc;
	reg error;

	//Temporary
	reg [3:0] register;

	// Instantiate the Unit Under Test (UUT)
	ld_st_shift_nbit uut (
		.clk(clk), 
		.clr(clr), 
		.set(set), 
		.ctrl(ctrl), 
		.ls(ls), 
		.rs(rs), 
		.reg_in(reg_in), 
		.reg_out(reg_out)
	);

	initial begin
		clk = 0;
		clr = 1;
		set = 1;
		reg_in = 0;
		ctrl = 0;
		ls = 0;
		rs = 0;
	end
	
	always begin
		//Generate CLOCK signal
		// Wait 100 ns for global reset to finish
		#10 clk = ~clk;

	end
	
	always									
		begin: testVector_loop
		integer c;
		for(c=0;c<256;c=c+1)
		begin: cLoop			//Equations generated by perl script truth_to_equation.pl - equations need simplification eventually
			#20	clr <= ~((c[5]&c[4]&c[3]&c[2]&~c[1]&c[0])|(c[5]&c[4]&c[3]&~c[2]&c[1]&~c[0])|(c[5]&c[4]&c[3]&~c[2]&~c[1]&c[0])|(c[5]&~c[4]&c[3]&c[2]&c[1]&~c[0])|(c[5]&~c[4]&c[3]&c[2]&~c[1]&c[0])|(c[5]&~c[4]&~c[3]&c[2]&c[1]&~c[0])|(c[5]&~c[4]&~c[3]&c[2]&~c[1]&c[0])|(~c[5]&c[4]&c[3]&~c[2]&~c[1]&c[0])|(~c[5]&c[4]&c[3]&~c[2]&~c[1]&~c[0])|(~c[5]&c[4]&~c[3]&c[2]&~c[1]&~c[0])|(~c[5]&~c[4]&c[3]&~c[2]&c[1]&~c[0])|(~c[5]&~c[4]&c[3]&~c[2]&~c[1]&c[0])|(~c[5]&~c[4]&~c[3]&c[2]&~c[1]&c[0]));
					set <= ~((c[5]&c[4]&c[3]&c[2]&~c[1]&c[0])|(c[5]&c[4]&~c[3]&c[2]&c[1]&~c[0])|(c[5]&c[4]&~c[3]&c[2]&~c[1]&c[0])|(c[5]&~c[4]&c[3]&~c[2]&c[1]&~c[0])|(c[5]&~c[4]&c[3]&~c[2]&~c[1]&c[0])|(c[5]&~c[4]&~c[3]&c[2]&c[1]&~c[0])|(c[5]&~c[4]&~c[3]&c[2]&~c[1]&c[0])|(~c[5]&c[4]&c[3]&c[2]&~c[1]&c[0])|(~c[5]&c[4]&c[3]&c[2]&~c[1]&~c[0])|(~c[5]&c[4]&~c[3]&c[2]&~c[1]&~c[0])|(~c[5]&~c[4]&c[3]&c[2]&c[1]&c[0])|(~c[5]&~c[4]&c[3]&c[2]&c[1]&~c[0])|(~c[5]&~c[4]&~c[3]&c[2]&~c[1]&c[0]));
					ls <= ~c[4];
					rs <= c[4]; 
					ctrl[0] <= c[5];
					ctrl[1] <= c[6];
					reg_in <= c[7:4];
		end
		//#250 error=1; //Signal end of run
	end
	
	always@(posedge clk) begin
		if(clr==1'b0) begin reg_out_tc=4'b0000; end
		else if(set==1'b0) begin reg_out_tc=4'b1111; end
		else if(ctrl==2'b00) begin //Store - Output does not change
			if(reg_out_tc==4'b0000) begin reg_out_tc=4'b0000; end
			else if(reg_out_tc==4'b0001) begin reg_out_tc=4'b0001; end
			else if(reg_out_tc==4'b0010) begin reg_out_tc=4'b0010; end
			else if(reg_out_tc==4'b0011) begin reg_out_tc=4'b0011; end
			else if(reg_out_tc==4'b0100) begin reg_out_tc=4'b0100; end
			else if(reg_out_tc==4'b0101) begin reg_out_tc=4'b0101; end
			else if(reg_out_tc==4'b0110) begin reg_out_tc=4'b0110; end
			else if(reg_out_tc==4'b0111) begin reg_out_tc=4'b0111; end
			else if(reg_out_tc==4'b1000) begin reg_out_tc=4'b1000; end
			else if(reg_out_tc==4'b1001) begin reg_out_tc=4'b1001; end
			else if(reg_out_tc==4'b1010) begin reg_out_tc=4'b1010; end
			else if(reg_out_tc==4'b1011) begin reg_out_tc=4'b1011; end
			else if(reg_out_tc==4'b1100) begin reg_out_tc=4'b1100; end
			else if(reg_out_tc==4'b1101) begin reg_out_tc=4'b1101; end
			else if(reg_out_tc==4'b1110) begin reg_out_tc=4'b1110; end
			else if(reg_out_tc==4'b1111) begin reg_out_tc=4'b1111; end
		end	
		else if(ctrl==2'b01) begin //Load
			if(reg_in==4'b0000) begin reg_out_tc=4'b0000; end
			else if(reg_in==4'b0001) begin reg_out_tc=4'b0001; end
			else if(reg_in==4'b0010) begin reg_out_tc=4'b0010; end
			else if(reg_in==4'b0011) begin reg_out_tc=4'b0011; end
			else if(reg_in==4'b0100) begin reg_out_tc=4'b0100; end
			else if(reg_in==4'b0101) begin reg_out_tc=4'b0101; end
			else if(reg_in==4'b0110) begin reg_out_tc=4'b0110; end
			else if(reg_in==4'b0111) begin reg_out_tc=4'b0111; end
			else if(reg_in==4'b1000) begin reg_out_tc=4'b1000; end
			else if(reg_in==4'b1001) begin reg_out_tc=4'b1001; end
			else if(reg_in==4'b1010) begin reg_out_tc=4'b1010; end
			else if(reg_in==4'b1011) begin reg_out_tc=4'b1011; end
			else if(reg_in==4'b1100) begin reg_out_tc=4'b1100; end
			else if(reg_in==4'b1101) begin reg_out_tc=4'b1101; end
			else if(reg_in==4'b1110) begin reg_out_tc=4'b1110; end
			else if(reg_in==4'b1111) begin reg_out_tc=4'b1111; end
		end	
		else if(ctrl==2'b10) begin //left shift
			if(ls==1'b1) begin
				if(reg_out_tc==4'b0000) begin reg_out_tc=4'b0001; end
				else if(reg_out_tc==4'b0001) begin reg_out_tc=4'b0011; end
				else if(reg_out_tc==4'b0010) begin reg_out_tc=4'b0101; end
				else if(reg_out_tc==4'b0011) begin reg_out_tc=4'b0111; end
				else if(reg_out_tc==4'b0100) begin reg_out_tc=4'b1001; end
				else if(reg_out_tc==4'b0101) begin reg_out_tc=4'b1011; end
				else if(reg_out_tc==4'b0110) begin reg_out_tc=4'b1101; end
				else if(reg_out_tc==4'b0111) begin reg_out_tc=4'b1111; end
				else if(reg_out_tc==4'b1000) begin reg_out_tc=4'b0001; end
				else if(reg_out_tc==4'b1001) begin reg_out_tc=4'b0011; end
				else if(reg_out_tc==4'b1010) begin reg_out_tc=4'b0101; end
				else if(reg_out_tc==4'b1011) begin reg_out_tc=4'b0111; end
				else if(reg_out_tc==4'b1100) begin reg_out_tc=4'b1001; end
				else if(reg_out_tc==4'b1101) begin reg_out_tc=4'b1011; end
				else if(reg_out_tc==4'b1110) begin reg_out_tc=4'b1101; end
				else if(reg_out_tc==4'b1111) begin reg_out_tc=4'b1111; end
			end
			else if(ls==1'b0) begin
				if(reg_out_tc==4'b0000) begin reg_out_tc=4'b0000; end
				else if(reg_out_tc==4'b0001) begin reg_out_tc=4'b0010; end
				else if(reg_out_tc==4'b0010) begin reg_out_tc=4'b0100; end
				else if(reg_out_tc==4'b0011) begin reg_out_tc=4'b0110; end
				else if(reg_out_tc==4'b0100) begin reg_out_tc=4'b1000; end
				else if(reg_out_tc==4'b0101) begin reg_out_tc=4'b1010; end
				else if(reg_out_tc==4'b0110) begin reg_out_tc=4'b1100; end
				else if(reg_out_tc==4'b0111) begin reg_out_tc=4'b1110; end
				else if(reg_out_tc==4'b1000) begin reg_out_tc=4'b0000; end
				else if(reg_out_tc==4'b1001) begin reg_out_tc=4'b0010; end
				else if(reg_out_tc==4'b1010) begin reg_out_tc=4'b0100; end
				else if(reg_out_tc==4'b1011) begin reg_out_tc=4'b0110; end
				else if(reg_out_tc==4'b1100) begin reg_out_tc=4'b1000; end
				else if(reg_out_tc==4'b1101) begin reg_out_tc=4'b1010; end
				else if(reg_out_tc==4'b1110) begin reg_out_tc=4'b1100; end
				else if(reg_out_tc==4'b1111) begin reg_out_tc=4'b1110; end
			end
		end
		else if(ctrl==2'b11) begin //Right Shift
			if(rs==2'b1) begin
				if(reg_out_tc==4'b0000) begin reg_out_tc=4'b1000; end
				else if(reg_out_tc==4'b0001) begin reg_out_tc=4'b1000; end
				else if(reg_out_tc==4'b0010) begin reg_out_tc=4'b1001; end
				else if(reg_out_tc==4'b0011) begin reg_out_tc=4'b1001; end
				else if(reg_out_tc==4'b0100) begin reg_out_tc=4'b1010; end
				else if(reg_out_tc==4'b0101) begin reg_out_tc=4'b1010; end
				else if(reg_out_tc==4'b0110) begin reg_out_tc=4'b1011; end
				else if(reg_out_tc==4'b0111) begin reg_out_tc=4'b1011; end
				else if(reg_out_tc==4'b1000) begin reg_out_tc=4'b1100; end
				else if(reg_out_tc==4'b1001) begin reg_out_tc=4'b1100; end
				else if(reg_out_tc==4'b1010) begin reg_out_tc=4'b1101; end
				else if(reg_out_tc==4'b1011) begin reg_out_tc=4'b1101; end
				else if(reg_out_tc==4'b1100) begin reg_out_tc=4'b1110; end
				else if(reg_out_tc==4'b1101) begin reg_out_tc=4'b1110; end
				else if(reg_out_tc==4'b1110) begin reg_out_tc=4'b1111; end
				else if(reg_out_tc==4'b1111) begin reg_out_tc=4'b1111; end
			end
			else if(rs==2'b0) begin
				if(reg_out_tc==4'b0000) begin reg_out_tc=4'b0000; end
				else if(reg_out_tc==4'b0001) begin reg_out_tc=4'b0000; end
				else if(reg_out_tc==4'b0010) begin reg_out_tc=4'b0001; end
				else if(reg_out_tc==4'b0011) begin reg_out_tc=4'b0001; end
				else if(reg_out_tc==4'b0100) begin reg_out_tc=4'b0010; end
				else if(reg_out_tc==4'b0101) begin reg_out_tc=4'b0010; end
				else if(reg_out_tc==4'b0110) begin reg_out_tc=4'b0011; end
				else if(reg_out_tc==4'b0111) begin reg_out_tc=4'b0011; end
				else if(reg_out_tc==4'b1000) begin reg_out_tc=4'b0100; end
				else if(reg_out_tc==4'b1001) begin reg_out_tc=4'b0100; end
				else if(reg_out_tc==4'b1010) begin reg_out_tc=4'b0101; end
				else if(reg_out_tc==4'b1011) begin reg_out_tc=4'b0101; end
				else if(reg_out_tc==4'b1100) begin reg_out_tc=4'b0110; end
				else if(reg_out_tc==4'b1101) begin reg_out_tc=4'b0110; end
				else if(reg_out_tc==4'b1110) begin reg_out_tc=4'b0111; end
				else if(reg_out_tc==4'b1111) begin reg_out_tc=4'b0111; end
			end
		end
		
		# 2 if(reg_out_tc == reg_out) begin error=0; end
		else  begin error=1; end
	end
      
endmodule

