library verilog;
use verilog.vl_types.all;
entity one_hot_fsm_vtf is
end one_hot_fsm_vtf;
