library verilog;
use verilog.vl_types.all;
entity mhvpis_vtf is
end mhvpis_vtf;
