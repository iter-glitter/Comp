library verilog;
use verilog.vl_types.all;
entity alu_nbit_vtf is
end alu_nbit_vtf;
