library verilog;
use verilog.vl_types.all;
entity alu_bitslice_vtf is
end alu_bitslice_vtf;
