`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    18:47:24 04/04/2013 
// Design Name: 
// Module Name:    processor 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module processor();



//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////// STAGE ONE ///////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
	
	
	
	
	
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////// STAGE TWO ///////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////	
	
	
endmodule
