library verilog;
use verilog.vl_types.all;
entity ls_reg_vtf is
end ls_reg_vtf;
